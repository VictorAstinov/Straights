-1203807219
h
79
8S 

h
79


h
79


c
80





6S 7S 
0
0
80
7S
0 1 2 3 4 5 6 7 8 9 10 11 12 13 
2
1
